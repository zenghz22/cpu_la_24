module csr_strl (
//output
        csr_re,
        csr_we,

//input
        op,
        exception,
        ecode);
    
endmodule